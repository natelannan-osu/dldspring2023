module sub (input logic [7:0] a, b, output logic [7:0] sum);

   assign sum = a - b;

endmodule // sub

